library verilog;
use verilog.vl_types.all;
entity TopDE_vlg_check_tst is
    port(
        AUD_ADCLRCK     : in     vl_logic;
        AUD_BCLK        : in     vl_logic;
        AUD_DACLRCK     : in     vl_logic;
        I2C_SDAT        : in     vl_logic;
        LCD_D           : in     vl_logic_vector(7 downto 0);
        OCLK            : in     vl_logic;
        OCLK100         : in     vl_logic;
        OCLK200         : in     vl_logic;
        OControlState   : in     vl_logic_vector(6 downto 0);
        ODAddress       : in     vl_logic_vector(31 downto 0);
        ODByteEnable    : in     vl_logic_vector(3 downto 0);
        ODReadData      : in     vl_logic_vector(31 downto 0);
        ODReadEnable    : in     vl_logic;
        ODWriteData     : in     vl_logic_vector(31 downto 0);
        ODWriteEnable   : in     vl_logic;
        OIAddress       : in     vl_logic_vector(31 downto 0);
        OIReadData      : in     vl_logic_vector(31 downto 0);
        OflagBank       : in     vl_logic_vector(7 downto 0);
        OwInstr         : in     vl_logic_vector(31 downto 0);
        OwPC            : in     vl_logic_vector(31 downto 0);
        OwRegDisp       : in     vl_logic_vector(31 downto 0);
        OwRegDispFPU    : in     vl_logic_vector(31 downto 0);
        OwRegDispSelect : in     vl_logic_vector(4 downto 0);
        PS2_KBCLK       : in     vl_logic;
        PS2_KBDAT       : in     vl_logic;
        SD_CMD          : in     vl_logic;
        SD_DAT          : in     vl_logic;
        SD_DAT3         : in     vl_logic;
        SRAM_DQ         : in     vl_logic_vector(31 downto 0);
        oAUD_DACDAT     : in     vl_logic;
        oAUD_XCK        : in     vl_logic;
        oHEX0_D         : in     vl_logic_vector(6 downto 0);
        oHEX0_DP        : in     vl_logic;
        oHEX1_D         : in     vl_logic_vector(6 downto 0);
        oHEX1_DP        : in     vl_logic;
        oHEX2_D         : in     vl_logic_vector(6 downto 0);
        oHEX2_DP        : in     vl_logic;
        oHEX3_D         : in     vl_logic_vector(6 downto 0);
        oHEX3_DP        : in     vl_logic;
        oHEX4_D         : in     vl_logic_vector(6 downto 0);
        oHEX4_DP        : in     vl_logic;
        oHEX5_D         : in     vl_logic_vector(6 downto 0);
        oHEX5_DP        : in     vl_logic;
        oHEX6_D         : in     vl_logic_vector(6 downto 0);
        oHEX6_DP        : in     vl_logic;
        oHEX7_D         : in     vl_logic_vector(6 downto 0);
        oHEX7_DP        : in     vl_logic;
        oI2C_SCLK       : in     vl_logic;
        oIRDA_TXD       : in     vl_logic;
        oLCD_BLON       : in     vl_logic;
        oLCD_EN         : in     vl_logic;
        oLCD_ON         : in     vl_logic;
        oLCD_RS         : in     vl_logic;
        oLCD_RW         : in     vl_logic;
        oLEDG           : in     vl_logic_vector(8 downto 0);
        oLEDR           : in     vl_logic_vector(17 downto 0);
        oSD_CLK         : in     vl_logic;
        oSRAM_A         : in     vl_logic_vector(18 downto 0);
        oSRAM_ADSC_N    : in     vl_logic;
        oSRAM_ADSP_N    : in     vl_logic;
        oSRAM_ADV_N     : in     vl_logic;
        oSRAM_BE_N      : in     vl_logic_vector(3 downto 0);
        oSRAM_CE1_N     : in     vl_logic;
        oSRAM_CE2       : in     vl_logic;
        oSRAM_CE3_N     : in     vl_logic;
        oSRAM_CLK       : in     vl_logic;
        oSRAM_GW_N      : in     vl_logic;
        oSRAM_OE_N      : in     vl_logic;
        oSRAM_WE_N      : in     vl_logic;
        oTD1_RESET_N    : in     vl_logic;
        oUART_CTS       : in     vl_logic;
        oUART_TXD       : in     vl_logic;
        oVGA_B          : in     vl_logic_vector(9 downto 0);
        oVGA_BLANK_N    : in     vl_logic;
        oVGA_CLOCK      : in     vl_logic;
        oVGA_G          : in     vl_logic_vector(9 downto 0);
        oVGA_HS         : in     vl_logic;
        oVGA_R          : in     vl_logic_vector(9 downto 0);
        oVGA_SYNC_N     : in     vl_logic;
        oVGA_VS         : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end TopDE_vlg_check_tst;
