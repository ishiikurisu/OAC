library verilog;
use verilog.vl_types.all;
entity TopDE_vlg_vec_tst is
end TopDE_vlg_vec_tst;
