library verilog;
use verilog.vl_types.all;
entity TopDE is
    port(
        altera_reserved_tms: in     vl_logic;
        altera_reserved_tck: in     vl_logic;
        altera_reserved_tdi: in     vl_logic;
        altera_reserved_tdo: out    vl_logic;
        iCLK_50         : in     vl_logic;
        iCLK_28         : in     vl_logic;
        iCLK_50_4       : in     vl_logic;
        iCLK_50_2       : in     vl_logic;
        iKEY            : in     vl_logic_vector(3 downto 0);
        iSW             : in     vl_logic_vector(17 downto 0);
        oLEDG           : out    vl_logic_vector(8 downto 0);
        oLEDR           : out    vl_logic_vector(17 downto 0);
        oHEX0_D         : out    vl_logic_vector(6 downto 0);
        oHEX1_D         : out    vl_logic_vector(6 downto 0);
        oHEX2_D         : out    vl_logic_vector(6 downto 0);
        oHEX3_D         : out    vl_logic_vector(6 downto 0);
        oHEX4_D         : out    vl_logic_vector(6 downto 0);
        oHEX5_D         : out    vl_logic_vector(6 downto 0);
        oHEX6_D         : out    vl_logic_vector(6 downto 0);
        oHEX7_D         : out    vl_logic_vector(6 downto 0);
        oHEX0_DP        : out    vl_logic;
        oHEX1_DP        : out    vl_logic;
        oHEX2_DP        : out    vl_logic;
        oHEX3_DP        : out    vl_logic;
        oHEX4_DP        : out    vl_logic;
        oHEX5_DP        : out    vl_logic;
        oHEX6_DP        : out    vl_logic;
        oHEX7_DP        : out    vl_logic;
        oVGA_CLOCK      : out    vl_logic;
        oVGA_HS         : out    vl_logic;
        oVGA_VS         : out    vl_logic;
        oVGA_BLANK_N    : out    vl_logic;
        oVGA_SYNC_N     : out    vl_logic;
        oVGA_R          : out    vl_logic_vector(9 downto 0);
        oVGA_G          : out    vl_logic_vector(9 downto 0);
        oVGA_B          : out    vl_logic_vector(9 downto 0);
        oTD1_RESET_N    : out    vl_logic;
        I2C_SDAT        : inout  vl_logic;
        oI2C_SCLK       : out    vl_logic;
        AUD_ADCLRCK     : inout  vl_logic;
        iAUD_ADCDAT     : in     vl_logic;
        AUD_DACLRCK     : out    vl_logic;
        oAUD_DACDAT     : out    vl_logic;
        AUD_BCLK        : inout  vl_logic;
        oAUD_XCK        : out    vl_logic;
        PS2_KBCLK       : inout  vl_logic;
        PS2_KBDAT       : inout  vl_logic;
        LCD_D           : inout  vl_logic_vector(7 downto 0);
        oLCD_ON         : out    vl_logic;
        oLCD_BLON       : out    vl_logic;
        oLCD_RW         : out    vl_logic;
        oLCD_EN         : out    vl_logic;
        oLCD_RS         : out    vl_logic;
        SRAM_DQ         : inout  vl_logic_vector(31 downto 0);
        oSRAM_A         : out    vl_logic_vector(18 downto 0);
        oSRAM_ADSC_N    : out    vl_logic;
        oSRAM_ADSP_N    : out    vl_logic;
        oSRAM_ADV_N     : out    vl_logic;
        oSRAM_BE_N      : out    vl_logic_vector(3 downto 0);
        oSRAM_CE1_N     : out    vl_logic;
        oSRAM_CE2       : out    vl_logic;
        oSRAM_CE3_N     : out    vl_logic;
        oSRAM_CLK       : out    vl_logic;
        oSRAM_GW_N      : out    vl_logic;
        oSRAM_OE_N      : out    vl_logic;
        oSRAM_WE_N      : out    vl_logic;
        oUART_TXD       : out    vl_logic;
        iUART_RXD       : in     vl_logic;
        oUART_CTS       : out    vl_logic;
        iUART_RTS       : in     vl_logic;
        oIRDA_TXD       : out    vl_logic;
        iIRDA_RXD       : in     vl_logic;
        OCLK            : out    vl_logic;
        OCLK100         : out    vl_logic;
        OCLK200         : out    vl_logic;
        OwRegDispSelect : out    vl_logic_vector(4 downto 0);
        OwPC            : out    vl_logic_vector(31 downto 0);
        OwInstr         : out    vl_logic_vector(31 downto 0);
        OwRegDisp       : out    vl_logic_vector(31 downto 0);
        OwRegDispFPU    : out    vl_logic_vector(31 downto 0);
        OflagBank       : out    vl_logic_vector(7 downto 0);
        ODReadEnable    : out    vl_logic;
        ODWriteEnable   : out    vl_logic;
        ODAddress       : out    vl_logic_vector(31 downto 0);
        ODWriteData     : out    vl_logic_vector(31 downto 0);
        ODReadData      : out    vl_logic_vector(31 downto 0);
        ODByteEnable    : out    vl_logic_vector(3 downto 0);
        OIAddress       : out    vl_logic_vector(31 downto 0);
        OIReadData      : out    vl_logic_vector(31 downto 0);
        OControlState   : out    vl_logic_vector(6 downto 0);
        SD_DAT3         : inout  vl_logic;
        SD_DAT          : inout  vl_logic;
        SD_CMD          : inout  vl_logic;
        oSD_CLK         : out    vl_logic
    );
end TopDE;
