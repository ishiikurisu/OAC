X <= A when S = '1' else B;