library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity ControlUnit is
	generic (
		WSIZE: natural := 32
	);
	port (
		
	);
end ControlUnit;

architecture rtl of ControlUnit is
	begin
	working: process()
	begin
		-- TODO Implement me!
	end process;
end rtl;
